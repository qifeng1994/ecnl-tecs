signature sOpenCloseSensor {
    void setDegreeOfOpeningDetectionStatus2_Yes( );
    void setDegreeOfOpeningDetectionStatus2_No( );
};
