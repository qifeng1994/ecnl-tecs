signature sLightingSystem {
    void setSceneControlSetting( );
    void getSceneControlSetting( );
    void getNumberThatCanAssignSceneControlSetting( );
};
