signature sGasLeakSensor {
    void getGasLeakOccurrenceStatus_Yes( );
    void getGasLeakOccurrenceStatus_No( );
};
