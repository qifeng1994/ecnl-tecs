signature sAirPollution {
    void setAirPollutionDetectionStatus_Yes( );
    void setAirPollutionDetectionStatus_No( );
};
