signature sDifferentialPressureSensor {
    void setMeasuredValueOfDifferentialPressure( );
};
