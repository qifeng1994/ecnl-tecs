signature sHouseholdSolarPowerGeneration {
    void setFitContractType_Fit( );
    void setFitContractType_NonFit( );
    void setFitContractType_NoSetting( );
    void getFitContractType_Fit( );
    void getFitContractType_NonFit( );
    void getFitContractType_NoSetting( );
    void getSelfConsumptionType_WithSelfConsumption( );
    void getSelfConsumptionType_WithoutSelfConsumption( );
    void getSelfConsumptionType_Unknown( );
    void getOutputPowerRestraintStatus_OngoingRestraint(outputPowerControl)( );
    void getOutputPowerRestraintStatus_OngoingRestraint(exceptOutputPowerControl)( );
    void getOutputPowerRestraintStatus_OngoingRestraint(reasonForRestraintIsUnknown)( );
    void getOutputPowerRestraintStatus_NotRestraining( );
    void getOutputPowerRestraintStatus_Unknown( );
    void getMeasuredInstantaneousAmountOfElectricityGenerated( );
    void getMeasuredCumulativeAmountOfElectricEnergyGenerated( );
};
