signature sGasHeatPumpTypeCommercialAirConditioner(outdoorUnit) {
};
