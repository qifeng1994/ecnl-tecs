signature sCombinationMicrowaveOven {
};
