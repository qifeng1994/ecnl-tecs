signature sBathroomHeaterAndDryer {
    void setBathroomDryerOperationSetting_Automatic( );
    void setBathroomDryerOperationSetting_Standard( );
    void getBathroomDryerOperationSetting_Automatic( );
    void getBathroomDryerOperationSetting_Standard( );
};
