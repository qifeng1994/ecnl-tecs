signature sDifferentialPressureSensor {
    void getMeasuredValueOfDifferentialPressure( );
};
