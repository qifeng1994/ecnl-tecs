signature sFuelCell {
    void getMeasuredInstantaneousPowerGenerationOutput( );
    void getMeasuredCumulativePowerGenerationOutput( );
    void setDesignatedPowerGenerationStatus_PowerGenerationAtTheMax.Rating( );
    void setDesignatedPowerGenerationStatus_LoadFollowingPowerGeneration( );
    void getDesignatedPowerGenerationStatus_PowerGenerationAtTheMax.Rating( );
    void getDesignatedPowerGenerationStatus_LoadFollowingPowerGeneration( );
};
