signature sRainSensor {
    void getRainDetectionStatus_Yes( );
    void getRainDetectionStatus_No( );
};
