signature sGasLeakSensor {
    void setGasLeakOccurrenceStatus_Yes( );
    void setGasLeakOccurrenceStatus_No( );
    void setGasLeakOccurrenceStatusResetting_Reset( );
};
