signature sMultipleInputPcs {
    void getSystemInterconnectedType_SystemInterconnectedType(reversePowerFlowAcceptable)( );
    void getSystemInterconnectedType_IndependentType( );
    void getSystemInterconnectedType_SystemInterconnectedType(reversePowerFlowNotAcceptable)( );
    void getMeasuredCumulativeAmountOfElectricEnergy(normalDirection)( );
    void getMeasuredCumulativeAmountOfElectricEnergy(reverseDirection)( );
    void getMeasuredInstantaneousElectricEnergy( );
};
