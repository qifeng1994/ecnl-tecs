signature sWaterFlowRate {
    void getFlowRate( );
};
