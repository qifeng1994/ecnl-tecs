signature sPowerDistributionBoard {
    void getMeasuredCumulativeAmountOfElectricEnergy(normalDirection)( );
    void getMeasuredCumulativeAmountOfElectricEnergy(reverseDirection)( );
};
