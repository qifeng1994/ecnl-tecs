signature sStorageBattery {
    void getAcEffectiveCapacity(charging)( );
    void getAcEffectiveCapacity(discharging)( );
    void getAcChargeableCapacity( );
    void getAcDischargeableCapacity( );
    void getAcChargeableElectricEnergy( );
    void getAcDischargeableElectricEnergy( );
    void getAcMeasuredCumulativeChargingElectricEnergy( );
    void getAcMeasuredCumulativeDischargingElectricEnergy( );
    void setAcChargeAmountSettingValue( );
    void getAcChargeAmountSettingValue( );
    void setAcDischargeAmountSettingValue( );
    void getAcDischargeAmountSettingValue( );
    void getChargingMethod_MaximumChargingElectricEnergyCharting( );
    void getChargingMethod_SurplusElectricEnergyCharging( );
    void getChargingMethod_DesignatedElectricEnergyCharging( );
    void getChargingMethod_DesignatedCurrentPowerCharging( );
    void getChargingMethod_Others( );
    void getDischargingMethod_MaximumDischargeElectricEnergyDischarging( );
    void getDischargingMethod_LoadFollowingDischarge( );
    void getDischargingMethod_DesignatedElectricEnergyDischarging( );
    void getDischargingMethod_DesignatedCurrentPowerDischarging( );
    void getDischargingMethod_Others( );
    void getBatteryType_Unknown( );
    void getBatteryType_Lead( );
    void getBatteryType_NiMh( );
    void getBatteryType_NiCd( );
    void getBatteryType_Lib( );
    void getBatteryType_Zinc( );
    void getBatteryType_Alkaline( );
};
