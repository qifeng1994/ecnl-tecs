signature sHighVoltageSmartElectricEnergyMeter {
    void getMonthlyMaximumElectricPowerDemand( );
    void getNumberOfEffectiveDigitsOfElectricPowerDemand( );
    void getCoefficient( );
    void getFixedDate( );
    void setDayForWhichTheHistoricalDataOfMeasuredCumulativeAmountsOfElectricEnergyIsToBeRetrieved( );
    void getDayForWhichTheHistoricalDataOfMeasuredCumulativeAmountsOfElectricEnergyIsToBeRetrieved( );
    void getNumberOfEffectiveDigitsForCumulativeAmountOfActiveElectricEnergy( );
};
