signature sAudio {
};
