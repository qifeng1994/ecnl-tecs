signature sBedPresenceSensor {
    void getBedPresenceDetectionStatus_Yes( );
    void getBedPresenceDetectionStatus_No( );
};
