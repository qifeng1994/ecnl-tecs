signature sSuperClass {
    void getOperationStatus_On( );
    void getOperationStatus_Off( );
    void getFaultStatus_Fault( );
    void getFaultStatus_NoFault( );
};
