signature sBathWaterLevelSensor {
    void getMeasuredValueOfBathWaterLevel( );
};
