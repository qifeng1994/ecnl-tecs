signature sElectricallyOperatedShade {
    void setOpenCloseSetting_Open( );
    void setOpenCloseSetting_Close( );
    void getOpenCloseSetting_Open( );
    void getOpenCloseSetting_Close( );
};
