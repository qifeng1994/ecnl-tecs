signature sMonoFunctionalLighting {
    void setIlluminanceLevel( );
};
