signature sElectricKey {
    void setLockSetting1_Lock( );
    void setLockSetting1_Unlock( );
    void getLockSetting1_Lock( );
    void getLockSetting1_Unlock( );
};
