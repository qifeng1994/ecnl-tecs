signature sVentilationFan {
};
