signature sCondensationSensor {
    void getCondensationDetectionStatus_Yes( );
    void getCondensationDetectionStatus_No( );
};
