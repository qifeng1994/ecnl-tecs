signature sGasSensor {
    void setGasDetectionStatus_Yes( );
    void setGasDetectionStatus_No( );
    void setMeasuredValueOfGasConcentration( );
};
