signature sPackageTypeCommercialAirConditioner(outdoorUnit) {
    void getMeasuredPowerConsumptionOfOutdoorUnit( );
    void getPossiblePowerSavingsForOutdoorUnits( );
    void setSettingsRestrictingPowerConsumptionOfOutdoorUnits( );
    void getSettingsRestrictingPowerConsumptionOfOutdoorUnits( );
};
