signature sWattHourMeter {
    void getCumulativeAmountsOfElectricEnergyMeasurementValue( );
};
