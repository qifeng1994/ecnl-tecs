signature sHumidifier {
};
