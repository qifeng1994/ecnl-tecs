signature sAirSpeedSensor {
    void getMeasuredValueOfAirSpeed( );
};
