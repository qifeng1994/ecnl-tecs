signature sFloorHeater {
};
