signature sExtendedLightingSystem {
    void setSceneControlSetting( );
    void getSceneControlSetting( );
    void getNumberThatCanAssignSceneControlSetting( );
    void getPowerConsumptionWhenFullyLighted( );
    void getPossiblePowerSavings( );
    void setPowerConsumptionLimitSetting( );
    void getPowerConsumptionLimitSetting( );
};
