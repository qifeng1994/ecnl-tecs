signature sInstantaneousWaterHeater {
    void getHotWaterHeatingStatus_Yes( );
    void getHotWaterHeatingStatus_No( );
    void getBathWaterHeaterStatus_Yes( );
    void getBathWaterHeaterStatus_No( );
    void setBathAutoModeSetting_On( );
    void setBathAutoModeSetting_Off( );
    void getBathAutoModeSetting_On( );
    void getBathAutoModeSetting_Off( );
};
