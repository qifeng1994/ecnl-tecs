signature sHumanDetectionSensor {
    void setHumanDetectionStatus_Yes( );
    void setHumanDetectionStatus_No( );
};
