signature sMonoFunctionalLighting {
};
