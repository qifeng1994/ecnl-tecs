signature sNetworkCamera {
    void setStillImagePhotographySetting_Shoot( );
};
