signature sWeightSensor {
    void getWeightDetectionStatus_Yes( );
    void getWeightDetectionStatus_No( );
};
