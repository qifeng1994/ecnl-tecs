signature sWaterLeakSensor {
    void getWaterLeakDetectionStatus_Yes( );
    void getWaterLeakDetectionStatus_No( );
};
