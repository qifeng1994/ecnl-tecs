signature sEvCharger {
    void setRatedChargeCapacity( );
    void setChargerDischargerType_AcCplt( );
    void setChargerDischargerType_AcHlcCharge( );
    void setChargerDischargerType_DcAaCharge( );
    void setChargerDischargerType_DcBbCharge( );
    void setChargerDischargerType_DcEeCharge( );
    void setChargerDischargerType_DcFfCharge( );
    void setVehicleConnectionConfirmation_ConnectionConfirmation( );
    void setChargeableCapacityOfVehicleMountedBattery( );
    void setRemainingChargeableCapacityOfVehicleMountedBattery( );
    void setUsedCapacityOfVehicleMountedBattery1( );
    void setRatedVoltage( );
    void setMeasuredInstantaneousChargingDischargingElectricEnergy( );
    void setMeasuredCumulativeAmountOfChargingElectricEnergy( );
    void setCumulativeAmountOfChargingElectricEnergyResetSetting_Reset( );
    void setOperationModeSetting_Charge( );
    void setOperationModeSetting_Standby( );
    void setOperationModeSetting_Idle( );
    void setOperationModeSetting_Other( );
    void setRemainingStoredElectricityOfVehicleMountedBattery1( );
    void setRemainingStoredElectricityOfVehicleMountedBattery3( );
    void setChargingAmountSetting( );
    void setChargingElectricEnergySetting( );
    void setChargingCurrentSetting( );
};
