signature sHumanBodyDetectionLocation1 {
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
        };
        
celltype tHumanBodyDetectionLocation1 {
        entry sHumanBodyDetectionLocation1 eHumanBodyDetectionLocation1;
        };
