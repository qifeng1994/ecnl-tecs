signature sMailingSensor {
    void getMailingDetectionStatus_Yes( );
    void getMailingDetectionStatus_No( );
};
