signature sWaterLevelSensor {
    void getMeasuredValueOfWaterLevel( );
};
