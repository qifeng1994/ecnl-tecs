signature sHybridWaterHeater {
    void setLinkageModeSettingForSolarPowerGeneration_ModeOff( );
    void setLinkageModeSettingForSolarPowerGeneration_HouseholdConsumption( );
    void setLinkageModeSettingForSolarPowerGeneration_PrioritizingElectricitySales( );
    void setLinkageModeSettingForSolarPowerGeneration_EconomicEfficiency( );
    void getLinkageModeSettingForSolarPowerGeneration_ModeOff( );
    void getLinkageModeSettingForSolarPowerGeneration_HouseholdConsumption( );
    void getLinkageModeSettingForSolarPowerGeneration_PrioritizingElectricitySales( );
    void getLinkageModeSettingForSolarPowerGeneration_EconomicEfficiency( );
};
