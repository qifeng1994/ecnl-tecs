signature sCrimePreventionSensor {
    void getInvasionOccurrenceStatus_Yes( );
    void getInvasionOccurrenceStatus_No( );
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
        };
        
celltype tCrimePreventionSensor {
        entry sCrimePreventionSensor eCrimePreventionSensor;
        };
