signature sIlluminanceSensor {
};
