signature sEvChargeAndDischargeSystem {
};
