signature sElectricEnergySensor {
    void getCumulativeAmountsOfElectricEnergy( );
};
