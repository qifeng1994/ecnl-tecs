signature sCigaretteSmokeSensor {
    void setSmoke(cigarette)DetectionStatus_Yes( );
    void setSmoke(cigarette)DetectionStatus_No( );
};
