signature sRainSensor {
    void setRainDetectionStatus_Yes( );
    void setRainDetectionStatus_No( );
};
