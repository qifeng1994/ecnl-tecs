signature sEngineCogeneration {
    void getMeasuredInstantaneousPowerGenerationOutput( );
    void getMeasuredCumulativePowerGenerationOutput( );
};
