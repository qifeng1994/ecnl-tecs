signature sLowVoltageSmartElectricEnergyMeter {
    void getNumberOfEffectiveDigitsForCumulativeAmountsOfElectricEnergy( );
    void getMeasuredCumulativeAmountOfElectricEnergy(normalDirection)( );
    void getMeasuredCumulativeAmountsOfElectricEnergy(reverseDirection)( );
    void setDayForWhichTheHistoricalDataOfMeasuredCumulativeAmountsOfElectricEnergyIsToBeRetrieved1( );
    void getDayForWhichTheHistoricalDataOfMeasuredCumulativeAmountsOfElectricEnergyIsToBeRetrieved1( );
    void getMeasuredInstantaneousElectricEnergy( );
};
