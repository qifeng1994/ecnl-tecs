signature sWaterOverflowSensor {
    void getWaterOverflowDetectionStatus_Yes( );
    void getWaterOverflowDetectionStatus_No( );
};
