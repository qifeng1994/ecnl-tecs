signature sRangeHood {
    void setVentilationAirFlowRateSetting_Automatic( );
    void setRangeHoodAutomaticSetting_Yes( );
    void setRangeHoodAutomaticSetting_No( );
    void setMeasuredValueOfIndoorTemperature( );
    void setMeasuredValueOfOutdoorTemperature( );
    void setMeasuredValueOfChargingAirTemperature( );
    void setMeasuredValueOfCookingTemperature( );
    void setMeasuredValueOfIndoorRelativeHumidity( );
    void setMeasuredValueOfOutdoorRelativeHumidity( );
    void setHumanDetectionStatus_Yes( );
    void setHumanDetectionStatus_No( );
    void setMeasuredValueOfCo2Concentration( );
    void setGasDetectionStatus_Yes( );
    void setGasDetectionStatus_No( );
    void setErrorDetectionMode_MotorError( );
    void setErrorDetectionMode_CurrentPlateDetection( );
    void setErrorDetectionMode_Normal( );
    void setErrorDetectionMode_Other( );
    void setLightingOperationSetting_Lighting( );
    void setLightingOperationSetting_LightsOut( );
    void setLightingOperationSetting_Flicker( );
    void setLightSourceColorSetting_IncandescentLampColor( );
    void setLightSourceColorSetting_White( );
    void setLightSourceColorSetting_DaylightWhite( );
    void setLightSourceColorSetting_DaylightColor( );
    void setLightSourceColorSetting_Other( );
    void setBrightnessLevelSetting( );
    void setLightingModeSetting_Automatic( );
    void setLightingModeSetting_NormalLighting( );
    void setLightingModeSetting_ColorLighting( );
};
