signature sAirCleaner {
};
