signature sGasHeatPumpTypeCommercialAirConditioner(indoorUnit) {
    void setThermoStatus_Yes( );
    void setThermoStatus_No( );
    void setOperationModeStatusDuringAutoOperation_Other( );
    void setOperationModeStatusDuringAutoOperation_Cooling( );
    void setOperationModeStatusDuringAutoOperation_Heating( );
    void setOperationModeStatusDuringAutoOperation_Dehumidification( );
    void setOperationModeStatusDuringAutoOperation_AirCirculation( );
    void setOperationModeSetting_Automatic( );
    void setOperationModeSetting_Cooling( );
    void setOperationModeSetting_Heating( );
    void setOperationModeSetting_Dehumidification( );
    void setOperationModeSetting_AirCirculation( );
    void setTemperatureSettingValue( );
    void setMeasuredTemperatureValueOfIndoorUnit( );
    void setPowerConsumptionRangeForIndoorUnits_Unknown( );
    void setPowerConsumptionRangeForIndoorUnits_LessThan50w( );
    void setPowerConsumptionRangeForIndoorUnits_50w100w( );
    void setPowerConsumptionRangeForIndoorUnits_100w150w( );
    void setPowerConsumptionRangeForIndoorUnits_150w200w( );
    void setPowerConsumptionRangeForIndoorUnits_EqualToOrMoreThan200w( );
};
