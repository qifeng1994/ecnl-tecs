signature sHumanBodyDetectionLocation1 {
};
