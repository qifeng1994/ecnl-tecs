signature sEmergencyButton {
    void getEmergencyOccurrenceStatus_Yes( );
    void getEmergencyOccurrenceStatus_No( );
};
