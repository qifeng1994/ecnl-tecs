signature sElectricallyOperatedBlindShade {
    void setOpenClose(extensionRetraction)Setting_Open( );
    void setOpenClose(extensionRetraction)Setting_Close( );
    void setOpenClose(extensionRetraction)Setting_Stop( );
    void getOpenClose(extensionRetraction)Setting_Open( );
    void getOpenClose(extensionRetraction)Setting_Close( );
    void getOpenClose(extensionRetraction)Setting_Stop( );
    void setDegreeOfOpeningLevel( );
    void getDegreeOfOpeningLevel( );
};
