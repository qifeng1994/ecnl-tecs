signature sSoundSensor {
    void setSoundDetectionStatus_Yes( );
    void setSoundDetectionStatus_No( );
    void setSoundDetectionHoldingTime( );
};
