signature sElectricLeakSensor {
    void getElectricLeakOccurrenceStatus_Yes( );
    void getElectricLeakOccurrenceStatus_No( );
};
