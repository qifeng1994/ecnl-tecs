signature sWaterFlowMeter {
    void getMeasuredCumulativeAmountOfFlowingWater( );
};
