signature sFlameSensor {
    void setFlameDetectionStatus_Yes( );
    void setFlameDetectionStatus_No( );
    void setFlameDetectionStatusResetting_Reset( );
};
