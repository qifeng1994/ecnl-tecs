signature sCurrentValueSensor {
    void setMeasuredCurrentValue1( );
    void setRatedVoltageToBeMeasured( );
    void setMeasuredCurrentValue2( );
};
