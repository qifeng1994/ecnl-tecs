signature sActivityAmountSensor {
};
