signature sCrimePreventionSensor {
    void getInvasionOccurrenceStatus_Yes( );
    void getInvasionOccurrenceStatus_No( );
};
