signature sBathroomHeaterAndDryer {
    void setOnTimerSetting1_On( );
    void setOnTimerSetting1_Off( );
    void setOffTimerSetting_On( );
    void setOffTimerSetting_Off( );
    void setVentilationOperationSetting_Automatic( );
    void setVentilationOperationSetting_Standard( );
    void setBathroomHeaterOperationSetting_Automatic( );
    void setBathroomHeaterOperationSetting_Standard( );
    void setBathroomDryerOperationSetting_Automatic( );
    void setBathroomDryerOperationSetting_Standard( );
    void setCoolAirCirculatorOperationSetting_Automatic( );
    void setCoolAirCirculatorOperationSetting_Standard( );
    void setMistSaunaOperationSetting_Automatic( );
    void setMistSaunaOperationSetting_Standard( );
    void setWaterMistOperationSetting_Automatic( );
    void setWaterMistOperationSetting_Standard( );
    void setMeasuredRelativeBathroomHumidity( );
    void setMeasuredBathroomTemperature( );
    void setVentilationAirFlowRateSetting_Automatic( );
    void setFilterCleaningReminderSignSetting_Lit( );
    void setFilterCleaningReminderSignSetting_NotLit( );
    void setHumanBodyDetectionStatus_Yes( );
    void setHumanBodyDetectionStatus_No( );
};
