signature sEarthquakeSensor {
    void getEarthquakeOccurrenceStatus_Yes( );
    void getEarthquakeOccurrenceStatus_No( );
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
};
celltype tEarthquakeSensor {
    entry sEarthquakeSensor eEarthquakeSensor;
};
