signature sSnowSensor {
    void getSnowDetectionStatus_Yes( );
    void getSnowDetectionStatus_No( );
};
