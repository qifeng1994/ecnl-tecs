signature sExtendedLightingSystem {
    void setIlluminanceLevelSetting( );
    void setSceneControlSetting( );
    void setNumberThatCanAssignSceneControlSetting( );
    void setPowerConsumptionWhenFullyLighted( );
    void setPossiblePowerSavings( );
    void setPowerConsumptionLimitSetting( );
    void setAutomaticOperationControllingSetting_On( );
    void setAutomaticOperationControllingSetting_Off( );
    void setFadingControlChangeTimeSetting( );
};
