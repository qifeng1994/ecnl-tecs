signature sVocSensor {
    void getMeasuredValueOfVocConcentration( );
};
