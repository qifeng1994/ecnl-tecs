signature sRefrigerator {
    void setQuickFreezeFunctionSetting_NormalOperation( );
    void setQuickFreezeFunctionSetting_QuickFreeze( );
    void setQuickFreezeFunctionSetting_StandbyForQuickFreezing( );
    void setQuickRefrigerationFunctionSetting_NormalOperation( );
    void setQuickRefrigerationFunctionSetting_QuickRefrigeration( );
    void setQuickRefrigerationFunctionSetting_StandbyForQuickRefrigeration( );
    void setIcemakerSetting_EnableIcemaker( );
    void setIcemakerSetting_DisableIcemaker( );
    void setIcemakerSetting_TemporarilyDisableIcemaker( );
    void setIcemakerOperationStatus_Yes( );
    void setIcemakerOperationStatus_No( );
    void setIcemakerTankStatus_WaterInTank( );
    void setIcemakerTankStatus_NoWater( );
    void setRefrigeratorCompartmentHumidificationFunctionSetting_On( );
    void setRefrigeratorCompartmentHumidificationFunctionSetting_Off( );
    void setVegetableCompartmentHumidificationFunctionSetting_On( );
    void setVegetableCompartmentHumidificationFunctionSetting_Off( );
    void setDeodorizationFunctionSetting_On( );
    void setDeodorizationFunctionSetting_Off( );
    void setDoorOpenCloseStatus_Open( );
    void setDoorOpenCloseStatus_Close( );
    void setDoorOpenWarning_Yes( );
    void setDoorOpenWarning_No( );
    void setRefrigeratorCompartmentDoorStatus_Open( );
    void setRefrigeratorCompartmentDoorStatus_Close( );
    void setFreezerCompartmentDoorStatus_Open( );
    void setFreezerCompartmentDoorStatus_Close( );
    void setIceCompartmentDoorStatus_Open( );
    void setIceCompartmentDoorStatus_Close( );
    void setVegetableCompartmentDoorStatus_Open( );
    void setVegetableCompartmentDoorStatus_Close( );
    void setMultiRefrigeratingModeCompartmentDoorStatus_Open( );
    void setMultiRefrigeratingModeCompartmentDoorStatus_Close( );
    void setMeasuredRefrigeratorCompartmentTemperature( );
    void setMeasuredFreezerCompartmentTemperature( );
    void setMeasuredSubzeroFreshCompartmentTemperature( );
    void setMeasuredVegetableCompartmentTemperature( );
    void setMeasuredMultiRefrigeratingModeCompartmentTemperature( );
    void setMeasuredElectricCurrentConsumption( );
    void setRatedPowerConsumption( );
    void setRefrigeratorCompartmentTemperatureSetting( );
    void setFreezerCompartmentTemperatureSetting( );
    void setIceTemperatureSetting( );
    void setVegetableCompartmentTemperatureSetting( );
    void setMultiRefrigeratingModeCompartmentTemperatureSetting( );
    void setRefrigeratorCompartmentTemperatureLevelSetting( );
    void setFreezerCompartmentTemperatureLevelSetting( );
    void setIceCompartmentTemperatureLevelSetting( );
    void setVegetableCompartmentTemperatureLevelSetting( );
    void setMultiRefrigeratingModeCompartmentTemperatureLevelSetting( );
};
