signature sOdorSensor {
    void getMeasuredOdorValue( );
};
