signature sSoundSensor {
    void getSoundDetectionStatus_Yes( );
    void getSoundDetectionStatus_No( );
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
        };
        
celltype tSoundSensor {
        entry sSoundSensor eSoundSensor;
        };
