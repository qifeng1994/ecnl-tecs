signature sBathWaterLevelSensor {
    void setBathWaterLevelOverDetectionThresholdLevel( );
    void setBathWaterLevelOverDetectionStatus_Yes( );
    void setBathWaterLevelOverDetectionStatus_No( );
    void setMeasuredValueOfBathWaterLevel( );
};
