signature sCookingHeater {
    void setAllStopSetting_StopAllHeating( );
};
