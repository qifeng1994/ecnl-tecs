signature sHouseholdSmallWindTurbinePowerGeneration {
    void getMeasuredInstantaneousAmountOfElectricityGenerated( );
    void getMeasuredCumulativeAmountOfElectricityGenerated( );
    void setBrakingStatus_On( );
    void setBrakingStatus_Off( );
    void getBrakingStatus_On( );
    void getBrakingStatus_Off( );
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
};
celltype tHouseholdSmallWindTurbinePowerGeneration {
    entry sHouseholdSmallWindTurbinePowerGeneration eHouseholdSmallWindTurbinePowerGeneration;
};
