signature sWeighingMachine {
};
