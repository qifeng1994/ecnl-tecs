signature sOxygenSensor {
    void getMeasuredValueOfOxygenConcentration( );
};
