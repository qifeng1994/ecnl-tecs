signature sTemperatureSensor {
    void setTemperatureValue( );
};
