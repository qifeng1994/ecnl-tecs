signature sSmartKerosenseMeter {
    void getMeasuredCumulativeKeroseneConsumption( );
};
