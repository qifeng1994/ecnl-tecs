signature sClothDryer {
};
