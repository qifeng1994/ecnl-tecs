signature sTelevision {
};
