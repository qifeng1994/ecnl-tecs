signature sBathroomHeaterAndDryer {
    void setBathroomDryerOperationSetting_Automatic( );
    void setBathroomDryerOperationSetting_Standard( );
    void getBathroomDryerOperationSetting_Automatic( );
    void getBathroomDryerOperationSetting_Standard( );
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
        };
        
celltype tBathroomHeaterAndDryer {
        entry sBathroomHeaterAndDryer eBathroomHeaterAndDryer;
        };
