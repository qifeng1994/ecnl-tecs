signature sRangeHood {
    void setVentilationAirFlowRateSetting_Automatic( );
    void getVentilationAirFlowRateSetting_Automatic( );
};
