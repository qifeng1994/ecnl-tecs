signature sHumanDetectionSensor {
    void getHumanDetectionStatus_Yes( );
    void getHumanDetectionStatus_No( );
};
