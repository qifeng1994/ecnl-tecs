signature sElectricHotWaterPot {
};
