signature sFlameSensor {
    void getFlameDetectionStatus_Yes( );
    void getFlameDetectionStatus_No( );
};
