signature sVocSensor {
    void setVocDetectionStatus_Yes( );
    void setVocDetectionStatus_No( );
    void setMeasuredValueOfVocConcentration( );
};
