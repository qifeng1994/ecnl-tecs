signature sCigaretteSmokeSensor {
    void getSmoke(cigarette)DetectionStatus_Yes( );
    void getSmoke(cigarette)DetectionStatus_No( );
};
