signature sGasMeter {
    void getCumulativeAmountOfGasConsumptionMeasurementValue( );
};
