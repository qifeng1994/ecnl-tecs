signature sController {
};
