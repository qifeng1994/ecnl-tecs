signature sIlluminanceSensor {
    void setIlluminanceValue1( );
    void setIlluminanceValue2( );
};
