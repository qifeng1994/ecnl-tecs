signature sCurrentValueSensor {
};
