signature sTemperatureSensor {
    void getTemperatureValue( );
};
