signature sCo2Sensor {
    void getMeasuredValueOfCo2Concentration( );
};
