signature sWattHourMeter {
    void setCumulativeAmountsOfElectricEnergyMeasurementValue( );
};
