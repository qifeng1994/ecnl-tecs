signature sBidetQuippedToilet(withElectricallyWarmedSeat) {
    void setHeaterSettingOfToiletSeat_On( );
    void setHeaterSettingOfToiletSeat_Off( );
    void getHeaterSettingOfToiletSeat_On( );
    void getHeaterSettingOfToiletSeat_Off( );
};
