signature sFanHeater {
    void setTemperatureSetValue( );
    void getTemperatureSetValue( );
};
