signature sVisitorSensor {
    void getVisitorDetectionStatus_Yes( );
    void getVisitorDetectionStatus_No( );
};
