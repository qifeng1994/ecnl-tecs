signature sDrEventController {
    void setNotificationIdDesignation( );
};
