signature sHumiditySensor {
    void getHumidityValue( );
};
