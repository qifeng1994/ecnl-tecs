signature sAirPollution {
    void getAirPollutionDetectionStatus_Yes( );
    void getAirPollutionDetectionStatus_No( );
};
