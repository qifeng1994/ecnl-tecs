signature sEarthquakeSensor {
    void getEarthquakeOccurrenceStatus_Yes( );
    void getEarthquakeOccurrenceStatus_No( );
};
