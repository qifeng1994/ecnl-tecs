signature sGardenSprinkler {
    void setSprinkleValveOpenCloseSetting_AutomaticOn( );
    void setSprinkleValveOpenCloseSetting_ManualOn( );
    void setSprinkleValveOpenCloseSetting_ManualOff( );
    void getSprinkleValveOpenCloseSetting_AutomaticOn( );
    void getSprinkleValveOpenCloseSetting_ManualOn( );
    void getSprinkleValveOpenCloseSetting_ManualOff( );
};
