signature sElectricallyOperatedShutter {
};
