signature sWeightSensor {
    void setWeightDetectionStatus_Yes( );
    void setWeightDetectionStatus_No( );
};
