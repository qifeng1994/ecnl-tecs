signature sOpenCloseSensor {
};
