signature sKerosenseMeter {
    void getMeasuredCumulativeAmountOfKeroseneConsumption( );
};
