signature sAirPressureSensor {
    void getAirPressureMeasurement( );
};
