signature sDishwasherAndDryer {
};
