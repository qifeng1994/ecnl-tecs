signature sRiceCooker {
    void setRiceCookingReservationSetting_On( );
    void setRiceCookingReservationSetting_Off( );
    void setCoverOpenCloseStatus_Open( );
    void setCoverOpenCloseStatus_Close( );
    void setRiceCookingStatus_Stop( );
    void setRiceCookingStatus_Preheating( );
    void setRiceCookingStatus_RiceCooking( );
    void setRiceCookingStatus_Steaming( );
