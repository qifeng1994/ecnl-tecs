signature sSnowSensor {
    void setSnowDetectionStatus_Yes( );
    void setSnowDetectionStatus_No( );
};
