signature sBidetQuippedToilet(withElectricallyWarmedSeat) {
    void setHeaterSettingOfToiletSeat_On( );
    void setHeaterSettingOfToiletSeat_Off( );
    void getHeaterSettingOfToiletSeat_On( );
    void getHeaterSettingOfToiletSeat_Off( );
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
        };
        
celltype tBidetQuippedToilet(withElectricallyWarmedSeat) {
        entry sBidetQuippedToilet(withElectricallyWarmedSeat) eBidetQuippedToilet(withElectricallyWarmedSeat);
        };
