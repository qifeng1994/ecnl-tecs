signature sCommercialShowCaseOutdoorUnit {
    void setOperationModeSetting_Cooling( );
    void setOperationModeSetting_NonCooling( );
};
