signature sElectricallyOperatedRainSlidingDoorShutter {
    void setOpenCloseSetting_Open( );
    void setOpenCloseSetting_Close( );
    void setOpenCloseSetting_Stop( );
    void getOpenCloseSetting_Open( );
    void getOpenCloseSetting_Close( );
    void getOpenCloseSetting_Stop( );
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
};
celltype tElectricallyOperatedRainSlidingDoorShutter {
    entry sElectricallyOperatedRainSlidingDoorShutter eElectricallyOperatedRainSlidingDoorShutter;
};
