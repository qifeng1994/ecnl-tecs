signature sElectricKey {
    void setLockSetting1_Lock( );
    void setLockSetting1_Unlock( );
    void getLockSetting1_Lock( );
    void getLockSetting1_Unlock( );
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
};
celltype tElectricKey {
    entry sElectricKey eElectricKey;
};
