signature sElectricallyOperatedWindow {
    void setTimerOperationSetting_On( );
    void setTimerOperationSetting_Off( );
    void setRegisteredTemperatureDetectionStatus_Yes( );
    void setRegisteredTemperatureDetectionStatus_No( );
    void setRainDetectionStatus_Yes( );
    void setRainDetectionStatus_No( );
    void setOpeningSpeedSetting_Low( );
    void setOpeningSpeedSetting_Middle( );
    void setOpeningSpeedSetting_High( );
    void setClosingSpeedSetting_Low( );
    void setClosingSpeedSetting_Middle( );
    void setClosingSpeedSetting_High( );
    void setOperationTime( );
    void setAutomaticOperationSetting_On( );
    void setAutomaticOperationSetting_Off( );
    void setOpenCloseSetting_Open( );
    void setOpenCloseSetting_Close( );
    void setOpenCloseSetting_Stop( );
    void setDegreeOfOpeningLevel( );
    void setOpeningClosingSpeedSetting_Low( );
    void setOpeningClosingSpeedSetting_Middle( );
    void setOpeningClosingSpeedSetting_High( );
    void setElectricLockSetting_Lock( );
    void setElectricLockSetting_Unlock( );
    void setRemoteOperationSettingStatus_On(permitted)( );
    void setRemoteOperationSettingStatus_Off(prohibited)( );
    void setSelectiveDegreeOfOpeningSetting_DegreeOfSettingPosition:Open( );
    void setSelectiveDegreeOfOpeningSetting_OperationTimeSettingValue:Open( );
    void setSelectiveDegreeOfOpeningSetting_OperationTimeSettingValue:Close( );
    void setSelectiveDegreeOfOpeningSetting_LocalSettingPosition( );
    void setOpenClosedStatus_FullyOpen( );
    void setOpenClosedStatus_FullyClosed( );
    void setOpenClosedStatus_Opening( );
    void setOpenClosedStatus_Closing( );
    void setOpenClosedStatus_StoppedHalfway( );
    void setOneTimeOpeningSpeedSetting_Low( );
    void setOneTimeOpeningSpeedSetting_Middle( );
    void setOneTimeOpeningSpeedSetting_High( );
    void setOneTimeOpeningSpeedSetting_None( );
    void setOneTimeClosingSpeedSetting_Low( );
    void setOneTimeClosingSpeedSetting_Middle( );
    void setOneTimeClosingSpeedSetting_High( );
    void setOneTimeClosingSpeedSetting_None( );
};
