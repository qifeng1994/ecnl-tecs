signature sFireSensor {
    void getFireOccurrenceDetectionStatus_Yes( );
    void getFireOccurrenceDetectionStatus_No( );
};
