signature sEvChargerAndDischarger {
    void getDischargeableCapacityOfVehicleMountedBattery1( );
    void getRemainingDischargeableCapacityOfVehicleMountedBattery1( );
    void getRemainingDischargeableCapacityOfVehicleMountedBattery3( );
    void getRatedChargeCapacity( );
    void getRatedDischargeCapacity( );
    void getChargerDischargerType_AcCplt( );
    void getChargerDischargerType_AcHlcCharge( );
    void getChargerDischargerType_AcHlcChargedischarge( );
    void getChargerDischargerType_DcAaCharge( );
    void getChargerDischargerType_DcAaChargedischarge( );
    void getChargerDischargerType_DcAaDischarge( );
    void getChargerDischargerType_DcBbCharge( );
    void getChargerDischargerType_DcBbChargedischarge( );
    void getChargerDischargerType_DcBbDischarge( );
    void getChargerDischargerType_DcEeCharge( );
    void getChargerDischargerType_DcEeChargedischarge( );
    void getChargerDischargerType_DcEeDischarge( );
    void getChargerDischargerType_DcFfCharge( );
    void getChargerDischargerType_DcFfChargedischarge( );
    void getChargerDischargerType_DcFfDischarge( );
    void setVehicleConnectionConfirmation_ConnectionConfirmation( );
    void getChargeableCapacityOfVehicleMountedBattery( );
    void getRemainingChargeableCapacityOfVehicleMountedBattery( );
    void getUsedCapacityOfVehicleMountedBattery1( );
    void getRemainingStoredElectricityOfVehicleMountedBattery1( );
    void getRemainingStoredElectricityOfVehicleMountedBattery3( );
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
};
celltype tEvChargerAndDischarger {
    entry sEvChargerAndDischarger eEvChargerAndDischarger;
};
