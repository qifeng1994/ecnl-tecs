signature sSoundSensor {
    void getSoundDetectionStatus_Yes( );
    void getSoundDetectionStatus_No( );
};
