signature sCallSensor {
    void getCallStatus_Yes( );
    void getCallStatus_No( );
};
