signature sBidetQuippedToilet(withElectricallyWarmedSeat) {
    void setHeaterSettingOfToiletSeat_On( );
    void setHeaterSettingOfToiletSeat_Off( );
    void setTemporalHaltSettingOfToiletSeat_Continuous( );
    void setTemporalHaltSettingOfToiletSeat_Once( );
    void setTemporalHaltSettingOfToiletSeat_NoSetting( );
    void setTemperatureLevelSettingOfRoomHeating_Low( );
    void setTemperatureLevelSettingOfRoomHeating_Medium( );
    void setTemperatureLevelSettingOfRoomHeating_High( );
    void setRoomHeatingSetting_On( );
    void setRoomHeatingSetting_Off( );
    void setRoomHeatingSetting_TimerMode( );
    void setRoomHeatingStatus_Yes( );
    void setRoomHeatingStatus_No( );
    void setSpecialOperationModeSetting_NoSetting( );
    void setSpecialOperationModeSetting_OverCoolPrevention( );
    void setHumanDetectionStatus_Yes( );
    void setHumanDetectionStatus_No( );
    void setSeatingDetectionStatus_Yes( );
    void setSeatingDetectionStatus_No( );
};
