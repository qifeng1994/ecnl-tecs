signature sAirPressureSensor {
    void setAirPressureMeasurement( );
};
