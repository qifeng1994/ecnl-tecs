signature sStorageBattery {
    void setAcEffectiveCapacity(charging)( );
    void setAcEffectiveCapacity(discharging)( );
    void setAcChargeableCapacity( );
    void setAcDischargeableCapacity( );
    void setAcChargeableElectricEnergy( );
    void setAcDischargeableElectricEnergy( );
    void setAcChargeUpperLimitSetting( );
    void setAcDischargeLowerLimitSetting( );
    void setAcMeasuredCumulativeChargingElectricEnergy( );
    void setAcMeasuredCumulativeDischargingElectricEnergy( );
    void setAcChargeAmountSettingValue( );
    void setAcDischargeAmountSettingValue( );
    void setChargingMethod_MaximumChargingElectricEnergyCharting( );
    void setChargingMethod_SurplusElectricEnergyCharging( );
    void setChargingMethod_DesignatedElectricEnergyCharging( );
    void setChargingMethod_DesignatedCurrentPowerCharging( );
    void setChargingMethod_Others( );
    void setDischargingMethod_MaximumDischargeElectricEnergyDischarging( );
    void setDischargingMethod_LoadFollowingDischarge( );
    void setDischargingMethod_DesignatedElectricEnergyDischarging( );
    void setDischargingMethod_DesignatedCurrentPowerDischarging( );
    void setDischargingMethod_Others( );
    void setAcRatedElectricEnergy( );
    void setReInterconnectionPermissionSetting_On( );
    void setReInterconnectionPermissionSetting_Off( );
    void setOperationPermissionSetting_On( );
    void setOperationPermissionSetting_Off( );
    void setIndependentOperationPermissionSetting_On( );
    void setIndependentOperationPermissionSetting_Off( );
    void setRatedElectricEnergy( );
    void setRatedCapacity( );
    void setRatedVoltage( );
    void setMeasuredInstantaneousChargingDischargingElectricEnergy( );
    void setMeasuredInstantaneousChargingDischargingCurrent( );
    void setMeasuredInstantaneousChargingDischargingVoltage( );
    void setMeasuredCumulativeDischargingElectricEnergy( );
    void setMeasuredCumulativeDischargingElectricEnergyResetSetting_Reset( );
    void setMeasuredCumulativeChargingElectricEnergy( );
    void setMeasuredCumulativeChargingElectricEnergyResetSetting_Reset( );
    void setChargingDischargingAmountSetting1( );
    void setChargingDischargingAmountSetting2( );
    void setRemainingStoredElectricity1( );
    void setRemainingStoredElectricity2( );
    void setRemainingStoredElectricity3( );
    void setBatteryStateOfHealth( );
    void setBatteryType_Unknown( );
    void setBatteryType_Lead( );
    void setBatteryType_NiMh( );
    void setBatteryType_NiCd( );
    void setBatteryType_Lib( );
    void setBatteryType_Zinc( );
    void setBatteryType_Alkaline( );
    void setChargingAmountSetting1( );
    void setDischargingAmountSetting1( );
    void setChargingAmountSetting2( );
    void setDischargingAmountSetting2( );
    void setChargingElectricEnergySetting( );
    void setDischargingElectricEnergySetting( );
    void setChargingCurrentSetting( );
    void setDischargingCurrentSetting( );
    void setRatedVoltage(independent)( );
};
