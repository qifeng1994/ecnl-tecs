signature sPackageTypeCommercialAirConditioner(outdoorUnit) {
    void setSpecialState_Yes( );
    void setSpecialState_No( );
    void setMeasuredOutdoorUnitTemperature( );
    void setMeasuredPowerConsumptionOfOutdoorUnit( );
    void setPossiblePowerSavingsForOutdoorUnits( );
    void setSettingsRestrictingPowerConsumptionOfOutdoorUnits( );
    void setMinimumPowerConsumptionForRestrictedOutdoorUnit( );
};
