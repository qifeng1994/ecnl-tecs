signature sBathHeatingStatusSensor {
    void getBathHeatingDetectionStatus_Yes( );
    void getBathHeatingDetectionStatus_No( );
};
