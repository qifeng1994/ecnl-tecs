signature sRefrigerator {
    void getDoorOpenCloseStatus_Open( );
    void getDoorOpenCloseStatus_Close( );
};
