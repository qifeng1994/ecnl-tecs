signature sElectricHeater {
    void setSetTemperatureValue( );
    void setSetTemperatureValue_Undefined( );
    void getSetTemperatureValue( );
    void getSetTemperatureValue_Undefined( );
};
