signature sGasSensor {
    void getMeasuredValueOfGasConcentration( );
};
