signature sDisplay {
};
