signature sNodeProfile {
    void getOperatingStatus_On( );
    void getOperatingStatus_Off( );
    void getNumberOfSelfNodeClasses( );
};
