signature sHotWaterHeatSourceEquipment {
};
