signature sKerosenseMeter {
    void setMeasuredCumulativeAmountOfKeroseneConsumption( );
};
