signature sParallelProcessingCombinationTypePowerControl {
};
