signature sWashingMachine {
};
