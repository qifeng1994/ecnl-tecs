signature sInstantaneousWaterHeater {
    void setOnTimerSetting_On( );
    void setOnTimerSetting_Off( );
    void setHotWaterHeatingStatus_Yes( );
    void setHotWaterHeatingStatus_No( );
    void setSetValueOfHotWaterTemperature( );
    void setHotWaterWarmerSetting_On( );
    void setHotWaterWarmerSetting_Off( );
    void setBathWaterVolumeSetting4( );
    void setBathWaterVolumeSetting4MaximumSettableLevel( );
    void setVolumeSetting( );
    void setMuteSetting_On( );
    void setMuteSetting_Off( );
    void setSetValueOfBathTemperature( );
    void setBathWaterHeaterStatus_Yes( );
    void setBathWaterHeaterStatus_No( );
    void setBathAutoModeSetting_On( );
    void setBathAutoModeSetting_Off( );
    void setBathAdditionalBoilUpOperationSetting_On( );
    void setBathAdditionalBoilUpOperationSetting_Off( );
    void setBathHotWaterAddingOperationSetting_On( );
    void setBathHotWaterAddingOperationSetting_Off( );
    void setBathWaterTemperatureLoweringOperationSetting_On( );
    void setBathWaterTemperatureLoweringOperationSetting_Off( );
    void setBathHotWaterVolumeSetting1( );
    void setShowerHotWaterSupplyStatus_Yes( );
    void setShowerHotWaterSupplyStatus_No( );
    void setKitchenHotWaterSupplyStatus_Yes( );
    void setKitchenHotWaterSupplyStatus_No( );
    void setHotWaterWarmerOnTimerReservationSetting_On( );
    void setHotWaterWarmerOnTimerReservationSetting_Off( );
    void setBathHotWaterVolumeSetting3( );
    void setBathOperationStatusMonitor_RunningHotWater( );
    void setBathOperationStatusMonitor_NoOperation( );
    void setBathOperationStatusMonitor_KeepingTemperature( );
};
