signature sElectricStorageHeater {
    void getHeatStorageOperationStatus_On( );
    void getHeatStorageOperationStatus_Off( );
    void setHeatStorageTemperatureSetting( );
    void getHeatStorageTemperatureSetting( );
    void getMeasuredStoredHeatTemperature( );
    void getMidnightPowerDurationSetting( );
    void setMidnightPowerStartTimeSetting( );
    void getMidnightPowerStartTimeSetting( );
    void getRadiationMethod_Yes( );
    void getRadiationMethod_No( );
};
