signature sFirstAidSensor {
    void setFirstAidOccurrenceStatus_Yes( );
    void setFirstAidOccurrenceStatus_No( );
    void setFirstAidOccurrenceStatusResetting_Reset( );
};
