signature sHouseholdSmallWindTurbinePowerGeneration {
    void getMeasuredInstantaneousAmountOfElectricityGenerated( );
    void getMeasuredCumulativeAmountOfElectricityGenerated( );
    void setBrakingStatus_On( );
    void setBrakingStatus_Off( );
    void getBrakingStatus_On( );
    void getBrakingStatus_Off( );
};
