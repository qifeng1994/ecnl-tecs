signature sFirstAidSensor {
    void getFirstAidOccurrenceStatus_Yes( );
    void getFirstAidOccurrenceStatus_No( );
};
