signature sMicromotionSensor {
    void getMicromotionDetectionStatus_Yes( );
    void getMicromotionDetectionStatus_No( );
};
