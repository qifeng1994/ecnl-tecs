signature sMultipleInputPcs {
    void getSystemInterconnectedType_SystemInterconnectedType(reversePowerFlowAcceptable)( );
    void getSystemInterconnectedType_IndependentType( );
    void getSystemInterconnectedType_SystemInterconnectedType(reversePowerFlowNotAcceptable)( );
    void getMeasuredCumulativeAmountOfElectricEnergy(normalDirection)( );
    void getMeasuredCumulativeAmountOfElectricEnergy(reverseDirection)( );
    void getMeasuredInstantaneousElectricEnergy( );
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
};
celltype tMultipleInputPcs {
    entry sMultipleInputPcs eMultipleInputPcs;
};
