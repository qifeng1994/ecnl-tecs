signature sSmartGasMeter {
};
