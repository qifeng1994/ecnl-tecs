signature sWasherAndDryer {
};
