signature sAirConditionerVentilationFan {
};
