signature sElectricWaterHeater {
    void getHotWaterSupplyStatus_Yes( );
    void getHotWaterSupplyStatus_No( );
    void setParticipationInEnergyShift_Participation( );
    void setParticipationInEnergyShift_NonParticipation( );
    void getParticipationInEnergyShift_Participation( );
    void getParticipationInEnergyShift_NonParticipation( );
    void getNumberOfEnergyShifts( );
    void setDaytimeHeatingShiftTime1( );
    void getDaytimeHeatingShiftTime1( );
    void setDaytimeHeatingShiftTime2( );
    void getDaytimeHeatingShiftTime2( );
    void setAutomaticBathWaterHeatingModeSetting_On( );
    void setAutomaticBathWaterHeatingModeSetting_Off( );
    void getAutomaticBathWaterHeatingModeSetting_On( );
    void getAutomaticBathWaterHeatingModeSetting_Off( );
};
