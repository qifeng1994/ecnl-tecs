signature sLpGasMeter {
};
