signature sGasMeter {
    void setCumulativeAmountOfGasConsumptionMeasurementValue( );
};
