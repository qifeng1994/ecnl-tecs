signature sBuzzar {
};
