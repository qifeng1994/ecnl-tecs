signature sGardenSprinkler {
    void setSprinkleValveOpenCloseSetting_AutomaticOn( );
    void setSprinkleValveOpenCloseSetting_ManualOn( );
    void setSprinkleValveOpenCloseSetting_ManualOff( );
    void getSprinkleValveOpenCloseSetting_AutomaticOn( );
    void getSprinkleValveOpenCloseSetting_ManualOn( );
    void getSprinkleValveOpenCloseSetting_ManualOff( );
    void setOperatingStatus_ON( );
    void getOperatingStatus_ON( );
    void setOperatingStatus_OFF( );
    void getOperatingStatus_OFF( );
    void setFaultStatus_Fault( );
    void getFaultStatus_Fault( );
    void setFaultStatus_NoFault( );
    void getFaultStatus_NoFault( );
        };
        
celltype tGardenSprinkler {
        entry sGardenSprinkler eGardenSprinkler;
        };
