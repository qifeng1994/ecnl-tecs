signature sLightingForSolidLightEmittingSource {
    void getNumberOfLightSources( );
};
