signature sWaterFlowRate {
    void setCumulativeFlowRate( );
    void setFlowRate( );
};
